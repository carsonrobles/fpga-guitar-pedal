`timescale 1ns / 1ps
`default_nettype none

module tri_wave_gen;


  //


endmodule
